library ieee;
use ieee.numeric_bit.all
