library ieee;
use ieee.std_logic_1164.all;

entity Exp8 is
  port(
    clock : in std_logic;
		Noturno, VeA, VeB, PdA, PdB				:	in std_logic; --Sinais externos (sensores ou comandos)
		reset								:	in std_logic; --Sinal de reset

    Q0, Q1, Q2  : out std_logic
  );
end entity;

architecture Exp8 of Exp8 is

  component CircuitoTemporizador is
    port(
      c1s, c5s, c1m : in std_logic;
      clock : in std_logic;

      cout  : out std_logic
    );
  end component;

  component FSMexp8 is
  	port(
  	--INPUTS
  		clock	:	in std_logic; --clocks para o circuito de 1 segundos, 5 segundos e 1 minuto
  		Noturno, VeA, VeB, PdA, PdB				:	in std_logic; --Sinais externos (sensores ou comandos)
  		reset								:	in std_logic; --Sinal de reset
  	--OUTPUTS
  		c1s, c5s, c1m:	out std_logic;
  		Q0, Q1, Q2	:	out std_logic
  		-- VmA, VdA, AmA					:	out std_logic; --Sinais de saida para semáforo A
  		-- VmB, VdB, AmB					:	out std_logic  --Sinais de saida para semaforo B
  	);
  end component;

  signal c1s, c5s, c1m  : std_logic;
  signal cout : std_logic;
  signal s0, s1, s2: std_logic;

begin

--  CT: CircuitoTemporizador port map(c1s => c1s, c5s => c5s, c1m => c1m, clock => clock, cout => cout);
--  FSM: FSMexp8 port map(clock => cout, Noturno => Noturno, VeA => VeA, VeB => VeB, PdA => PdA, PdB => PdB, reset => reset, c1s => c1s, c5s => c5s, c1m => c1m, Q0 => s0, Q1 => s1, Q2 => s2);


  CT: CircuitoTemporizador port map(c1s, c5s, c1m, clock, cout);
  FSM: FSMexp8 port map(cout, Noturno, VeA, VeB, PdA, PdB, reset, c1s, c5s, c1m, s0, s1, s2);


  Q0 <= s0;
  Q1 <= s1;
  Q2 <= s2;

end architecture;
